
`timescale 1ns / 1ps

module daddaTree (
  input logic [5:0][12:0] ops,
  output logic [18:0] result
);
  logic [5:0][17:0] M1;

  logic x;

  assign x = 1;


endmodule
